// Verilog
// c864
// Ninputs 72
// Noutputs 14
// NtotalGates 320
// NOT1 80
// NAND2 128
// NOR2 38
// AND9 6
// XOR2 36
// NAND4 28
// AND8 2
// NAND3 2

module c864 (N11,  N14,  N18,  N111, N114, N117, N121, N124, N127, N130,
             N134, N137, N140, N143, N147, N150, N153, N156, N160, N163,
             N166, N169, N173, N176, N179, N182, N186, N189, N192, N195,
             N199, N1102,N1105,N1108,N1112,N1115,N1223,N1329,N1370,N1421,
             N1430,N1431,N1432,
             N21,  N24,  N28,  N211, N214, N217, N221, N224, N227, N230,
             N234, N237, N240, N243, N247, N250, N253, N256, N260, N263,
             N266, N269, N273, N276, N279, N282, N286, N289, N292, N295,
             N299, N2102,N2105,N2108,N2112,N2115,N2223,N2329,N2370,N2421,
             N2430,N2431,N2432
);

input N11, N14,  N18,  N111, N114, N117, N121, N124, N127, N130,
      N134,N137, N140, N143, N147, N150, N153, N156, N160, N163,
      N166,N169, N173, N176, N179, N182, N186, N189, N192, N195,
      N199,N1102,N1105,N1108,N1112,N1115,
      N21, N24,  N28,  N211, N214, N217, N221, N224, N227, N230,
      N234,N237, N240, N243, N247, N250, N253, N256, N260, N263,
      N266,N269, N273, N276, N279, N282, N286, N289, N292, N295,
      N299,N2102,N2105,N2108,N2112,N2115;

output N1223,N1329,N1370,N1421,N1430,N1431,N1432,
       N2223,N2329,N2370,N2421,N2430,N2431,N2432;

wire N1118,N1119,N1122,N1123,N1126,N1127,N1130,N1131,N1134,N1135,
     N1138,N1139,N1142,N1143,N1146,N1147,N1150,N1151,N1154,N1157,
     N1158,N1159,N1162,N1165,N1168,N1171,N1174,N1177,N1180,N1183,
     N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,
     N1194,N1195,N1196,N1197,N1198,N1199,N1203,N1213,N1224,N1227,
     N1230,N1233,N1236,N1239,N1242,N1243,N1246,N1247,N1250,N1251,
     N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1263,N1264,N1267,
     N1270,N1273,N1276,N1279,N1282,N1285,N1288,N1289,N1290,N1291,
     N1292,N1293,N1294,N1295,N1296,N1300,N1301,N1302,N1303,N1304,
     N1305,N1306,N1307,N1308,N1309,N1319,N1330,N1331,N1332,N1333,
     N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,
     N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,
     N1354,N1355,N1356,N1357,N1360,N1371,N1372,N1373,N1374,N1375,
     N1376,N1377,N1378,N1379,N1380,N1381,N1386,N1393,N1399,N1404,
     N1407,N1411,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1422,
     N1425,N1428,N1429,
     N2118,N2119,N2122,N2123,N2126,N2127,N2130,N2131,N2134,N2135,
     N2138,N2139,N2142,N2143,N2146,N2147,N2150,N2151,N2154,N2157,
     N2158,N2159,N2162,N2165,N2168,N2171,N2174,N2177,N2180,N2183,
     N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,
     N2194,N2195,N2196,N2197,N2198,N2199,N2203,N2213,N2224,N2227,
     N2230,N2233,N2236,N2239,N2242,N2243,N2246,N2247,N2250,N2251,
     N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2263,N2264,N2267,
     N2270,N2273,N2276,N2279,N2282,N2285,N2288,N2289,N2290,N2291,
     N2292,N2293,N2294,N2295,N2296,N2300,N2301,N2302,N2303,N2304,
     N2305,N2306,N2307,N2308,N2309,N2319,N2330,N2331,N2332,N2333,
     N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,
     N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,
     N2354,N2355,N2356,N2357,N2360,N2371,N2372,N2373,N2374,N2375,
     N2376,N2377,N2378,N2379,N2380,N2381,N2386,N2393,N2399,N2404,
     N2407,N2411,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2422,
     N2425,N2428,N2429;

not  NOT1_11    (N1118, N11);
not  NOT1_12    (N1119, N14);
not  NOT1_13    (N1122, N111);
not  NOT1_14    (N1123, N117);
not  NOT1_15    (N1126, N124);
not  NOT1_16    (N1127, N130);
not  NOT1_17    (N1130, N137);
not  NOT1_18    (N1131, N143);
not  NOT1_19    (N1134, N150);	
not  NOT1_110   (N1135, N156);
not  NOT1_111   (N1138, N163);
not  NOT1_112   (N1139, N169);
not  NOT1_113   (N1142, N176);
not  NOT1_114   (N1143, N182);
not  NOT1_115   (N1146, N189);
not  NOT1_116   (N1147, N195);
not  NOT1_117   (N1150, N1102);
not  NOT1_118   (N1151, N1108);
not  NOT1_147   (N1203, N1199);
not  NOT1_148   (N1213, N1199);
not  NOT1_149   (N1223, N1199);
not  NOT1_187   (N1300, N1263);
not  NOT1_188   (N1301, N1288);
not  NOT1_189   (N1302, N1289);
not  NOT1_190   (N1303, N1290);
not  NOT1_191   (N1304, N1291);
not  NOT1_192   (N1305, N1292);
not  NOT1_193   (N1306, N1293);
not  NOT1_194   (N1307, N1294);
not  NOT1_195   (N1308, N1295);
not  NOT1_196   (N1309, N1296);
not  NOT1_197   (N1319, N1296);
not  NOT1_198   (N1329, N1296);
not  NOT1_1147  (N1415, N1380);
not  NOT1_1149  (N1417, N1393);
not  NOT1_1150  (N1418, N1404);
not  NOT1_1151  (N1419, N1407);
not  NOT1_1152  (N1420, N1411);
not  NOT1_1127  (N1360, N1357);
not  NOT1_1128  (N1370, N1357);
nor  NOR2_120   (N1157, N18,   N1119);
nor  NOR2_121   (N1158, N114,  N1119);
nor  NOR2_130   (N1183, N121,  N1123);
nor  NOR2_131   (N1184, N127,  N1123);
nor  NOR2_132   (N1185, N134,  N1127);
nor  NOR2_133   (N1186, N140,  N1127);
nor  NOR2_134   (N1187, N147,  N1131);
nor  NOR2_135   (N1188, N153,  N1131);
nor  NOR2_136   (N1189, N160,  N1135);
nor  NOR2_137   (N1190, N166,  N1135);
nor  NOR2_138   (N1191, N173,  N1139);
nor  NOR2_139   (N1192, N179,  N1139);
nor  NOR2_140   (N1193, N186,  N1143);
nor  NOR2_141   (N1194, N192,  N1143);
nor  NOR2_142   (N1195, N199,  N1147);
nor  NOR2_143   (N1196, N1105, N1147);
nor  NOR2_144   (N1197, N1112, N1151);
nor  NOR2_145   (N1198, N1115, N1151);
nor  NOR2_1153  (N1421, N1415, N1416);
xor  XOR2_150   (N1224, N1203, N1154);
xor  XOR2_151   (N1227, N1203, N1159);
xor  XOR2_152   (N1230, N1203, N1162);
xor  XOR2_153   (N1233, N1203, N1165);
xor  XOR2_154   (N1236, N1203, N1168);
xor  XOR2_155   (N1239, N1203, N1171);
xor  XOR2_157   (N1243, N1203, N1174);
xor  XOR2_159   (N1247, N1203, N1177);
xor  XOR2_161   (N1251, N1203, N1180);
xor  XOR2_199   (N1330, N1309, N1260);
xor  XOR2_1100  (N1331, N1309, N1264);
xor  XOR2_1101  (N1332, N1309, N1267);
xor  XOR2_1102  (N1333, N1309, N1270);
xor  XOR2_1104  (N1335, N1309, N1273);
xor  XOR2_1106  (N1337, N1309, N1276);
xor  XOR2_1108  (N1339, N1309, N1279);
xor  XOR2_1110  (N1341, N1309, N1282);
xor  XOR2_1112  (N1343, N1309, N1285);
nand NAND2_1103 (N1334, N18,   N1319);
nand NAND2_1105 (N1336, N1319, N121);
nand NAND2_1107 (N1338, N1319, N134);
nand NAND2_1109 (N1340, N1319, N147);
nand NAND2_1111 (N1342, N1319, N160);
nand NAND2_1154 (N1422, N1386, N1417);
nand NAND2_119  (N1154, N1118, N14);
nand NAND2_122  (N1159, N1122, N117);
nand NAND2_123  (N1162, N1126, N130);
nand NAND2_124  (N1165, N1130, N143);
nand NAND2_125  (N1168, N1134, N156);
nand NAND2_126  (N1171, N1138, N169);
nand NAND2_127  (N1174, N1142, N182);
nand NAND2_128  (N1177, N1146, N195);
nand NAND2_129  (N1180, N1150, N1108);
nand NAND2_156  (N1242, N11,   N1213);
nand NAND2_158  (N1246, N1213, N111);
nand NAND2_160  (N1250, N1213, N124);
nand NAND2_162  (N1254, N1213, N137);
nand NAND2_163  (N1255, N1213, N150);
nand NAND2_164  (N1256, N1213, N163);
nand NAND2_165  (N1257, N1213, N176);
nand NAND2_166  (N1258, N1213, N189);
nand NAND2_167  (N1259, N1213, N1102);
nand NAND2_168  (N1260, N1224, N1157);
nand NAND2_169  (N1263, N1224, N1158);
nand NAND2_170  (N1264, N1227, N1183);
nand NAND2_171  (N1267, N1230, N1185);
nand NAND2_172  (N1270, N1233, N1187);
nand NAND2_173  (N1273, N1236, N1189);
nand NAND2_174  (N1276, N1239, N1191);
nand NAND2_175  (N1279, N1243, N1193);
nand NAND2_176  (N1282, N1247, N1195);
nand NAND2_177  (N1285, N1251, N1197);
nand NAND2_178  (N1288, N1227, N1184);
nand NAND2_179  (N1289, N1230, N1186);
nand NAND2_180  (N1290, N1233, N1188);
nand NAND2_181  (N1291, N1236, N1190);
nand NAND2_182  (N1292, N1239, N1192);
nand NAND2_183  (N1293, N1243, N1194);
nand NAND2_184  (N1294, N1247, N1196);
nand NAND2_185  (N1295, N1251, N1198);
nand NAND2_1113 (N1344, N1319, N173);
nand NAND2_1114 (N1345, N1319, N186);
nand NAND2_1115 (N1346, N1319, N199);
nand NAND2_1116 (N1347, N1319, N1112);
nand NAND2_1117 (N1348, N1330, N1300);
nand NAND2_1118 (N1349, N1331, N1301);
nand NAND2_1119 (N1350, N1332, N1302);
nand NAND2_1120 (N1351, N1333, N1303);
nand NAND2_1121 (N1352, N1335, N1304);
nand NAND2_1122 (N1353, N1337, N1305);
nand NAND2_1123 (N1354, N1339, N1306);
nand NAND2_1124 (N1355, N1341, N1307);
nand NAND2_1125 (N1356, N1343, N1308);
nand NAND2_1129 (N1371, N114,  N1360);
nand NAND2_1130 (N1372, N1360, N127);
nand NAND2_1131 (N1373, N1360, N140);
nand NAND2_1132 (N1374, N1360, N153);
nand NAND2_1133 (N1375, N1360, N166);
nand NAND2_1134 (N1376, N1360, N179);
nand NAND2_1135 (N1377, N1360, N192);
nand NAND2_1136 (N1378, N1360, N1105);
nand NAND2_1137 (N1379, N1360, N1115);
nand NAND3_1156 (N1428, N1399, N1393, N1419);
nand NAND4_1138 (N1380, N14,   N1242, N1334, N1371);
nand NAND4_1139 (N1381, N1246, N1336, N1372, N117);
nand NAND4_1140 (N1386, N1250, N1338, N1373, N130);
nand NAND4_1141 (N1393, N1254, N1340, N1374, N143);
nand NAND4_1142 (N1399, N1255, N1342, N1375, N156);
nand NAND4_1143 (N1404, N1256, N1344, N1376, N169);
nand NAND4_1144 (N1407, N1257, N1345, N1377, N182);
nand NAND4_1145 (N1411, N1258, N1346, N1378, N195);
nand NAND4_1146 (N1414, N1259, N1347, N1379, N1108);
nand NAND4_1155 (N1425, N1386, N1393, N1418, N1399);
nand NAND4_1157 (N1429, N1386, N1393, N1407, N1420);
nand NAND4_1158 (N1430, N1381, N1386, N1422, N1399);
nand NAND4_1159 (N1431, N1381, N1386, N1425, N1428);
nand NAND4_1160 (N1432, N1381, N1422, N1425, N1429);
and  AND8_1148  (N1416, N1381, N1386, N1393, N1399, N1404, N1407, N1411, N1414);
and  AND9_146   (N1199, N1154, N1159, N1162, N1165, N1168, N1171, N1174, N1177, N1180);
and  AND9_186   (N1296, N1260, N1264, N1267, N1270, N1273, N1276, N1279, N1282, N1285);
and  AND9_1126  (N1357, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356);

not  NOT1_21    (N2118, N21);
not  NOT1_22    (N2119, N24);
not  NOT1_23    (N2122, N211);
not  NOT1_24    (N2123, N217);
not  NOT1_25    (N2126, N224);
not  NOT1_26    (N2127, N230);
not  NOT1_27    (N2130, N237);
not  NOT1_28    (N2131, N243);
not  NOT1_29    (N2134, N250);	
not  NOT1_210   (N2135, N256);
not  NOT1_211   (N2138, N263);
not  NOT1_212   (N2139, N269);
not  NOT1_213   (N2142, N276);
not  NOT1_214   (N2143, N282);
not  NOT1_215   (N2146, N289);
not  NOT1_216   (N2147, N295);
not  NOT1_217   (N2150, N2102);
not  NOT1_218   (N2151, N2108);
not  NOT1_247   (N2203, N2199);
not  NOT1_248   (N2213, N2199);
not  NOT1_249   (N2223, N2199);
not  NOT1_287   (N2300, N2263);
not  NOT1_288   (N2301, N2288);
not  NOT1_289   (N2302, N2289);
not  NOT1_290   (N2303, N2290);
not  NOT1_291   (N2304, N2291);
not  NOT1_292   (N2305, N2292);
not  NOT1_293   (N2306, N2293);
not  NOT1_294   (N2307, N2294);
not  NOT1_295   (N2308, N2295);
not  NOT1_296   (N2309, N2296);
not  NOT1_297   (N2319, N2296);
not  NOT1_298   (N2329, N2296);
not  NOT1_2147  (N2415, N2380);
not  NOT1_2149  (N2417, N2393);
not  NOT1_2150  (N2418, N2404);
not  NOT1_2151  (N2419, N2407);
not  NOT1_2152  (N2420, N2411);
not  NOT1_2127  (N2360, N2357);
not  NOT1_2128  (N2370, N2357);
nor  NOR2_220   (N2157, N28,   N2119);
nor  NOR2_221   (N2158, N214,  N2119);
nor  NOR2_230   (N2183, N221,  N2123);
nor  NOR2_231   (N2184, N227,  N2123);
nor  NOR2_232   (N2185, N234,  N2127);
nor  NOR2_233   (N2186, N240,  N2127);
nor  NOR2_234   (N2187, N247,  N2131);
nor  NOR2_235   (N2188, N253,  N2131);
nor  NOR2_236   (N2189, N260,  N2135);
nor  NOR2_237   (N2190, N266,  N2135);
nor  NOR2_238   (N2191, N273,  N2139);
nor  NOR2_239   (N2192, N279,  N2139);
nor  NOR2_240   (N2193, N286,  N2143);
nor  NOR2_241   (N2194, N292,  N2143);
nor  NOR2_242   (N2195, N299,  N2147);
nor  NOR2_243   (N2196, N2105, N2147);
nor  NOR2_244   (N2197, N2112, N2151);
nor  NOR2_245   (N2198, N2115, N2151);
nor  NOR2_2153  (N2421, N2415, N2416);
xor  XOR2_250   (N2224, N2203, N2154);
xor  XOR2_251   (N2227, N2203, N2159);
xor  XOR2_252   (N2230, N2203, N2162);
xor  XOR2_253   (N2233, N2203, N2165);
xor  XOR2_254   (N2236, N2203, N2168);
xor  XOR2_255   (N2239, N2203, N2171);
xor  XOR2_257   (N2243, N2203, N2174);
xor  XOR2_259   (N2247, N2203, N2177);
xor  XOR2_261   (N2251, N2203, N2180);
xor  XOR2_299   (N2330, N2309, N2260);
xor  XOR2_2100  (N2331, N2309, N2264);
xor  XOR2_2101  (N2332, N2309, N2267);
xor  XOR2_2102  (N2333, N2309, N2270);
xor  XOR2_2104  (N2335, N2309, N2273);
xor  XOR2_2106  (N2337, N2309, N2276);
xor  XOR2_2108  (N2339, N2309, N2279);
xor  XOR2_2110  (N2341, N2309, N2282);
xor  XOR2_2112  (N2343, N2309, N2285);
nand NAND2_2103 (N2334, N28,   N2319);
nand NAND2_2105 (N2336, N2319, N221);
nand NAND2_2107 (N2338, N2319, N234);
nand NAND2_2109 (N2340, N2319, N247);
nand NAND2_2111 (N2342, N2319, N260);
nand NAND2_2154 (N2422, N2386, N2417);
nand NAND2_219  (N2154, N2118, N24);
nand NAND2_222  (N2159, N2122, N217);
nand NAND2_223  (N2162, N2126, N230);
nand NAND2_224  (N2165, N2130, N243);
nand NAND2_225  (N2168, N2134, N256);
nand NAND2_226  (N2171, N2138, N269);
nand NAND2_227  (N2174, N2142, N282);
nand NAND2_228  (N2177, N2146, N295);
nand NAND2_229  (N2180, N2150, N2108);
nand NAND2_256  (N2242, N21,   N2213);
nand NAND2_258  (N2246, N2213, N211);
nand NAND2_260  (N2250, N2213, N224);
nand NAND2_262  (N2254, N2213, N237);
nand NAND2_263  (N2255, N2213, N250);
nand NAND2_264  (N2256, N2213, N263);
nand NAND2_265  (N2257, N2213, N276);
nand NAND2_266  (N2258, N2213, N289);
nand NAND2_267  (N2259, N2213, N2102);
nand NAND2_268  (N2260, N2224, N2157);
nand NAND2_269  (N2263, N2224, N2158);
nand NAND2_270  (N2264, N2227, N2183);
nand NAND2_271  (N2267, N2230, N2185);
nand NAND2_272  (N2270, N2233, N2187);
nand NAND2_273  (N2273, N2236, N2189);
nand NAND2_274  (N2276, N2239, N2191);
nand NAND2_275  (N2279, N2243, N2193);
nand NAND2_276  (N2282, N2247, N2195);
nand NAND2_277  (N2285, N2251, N2197);
nand NAND2_278  (N2288, N2227, N2184);
nand NAND2_279  (N2289, N2230, N2186);
nand NAND2_280  (N2290, N2233, N2188);
nand NAND2_281  (N2291, N2236, N2190);
nand NAND2_282  (N2292, N2239, N2192);
nand NAND2_283  (N2293, N2243, N2194);
nand NAND2_284  (N2294, N2247, N2196);
nand NAND2_285  (N2295, N2251, N2198);
nand NAND2_2113 (N2344, N2319, N273);
nand NAND2_2114 (N2345, N2319, N286);
nand NAND2_2115 (N2346, N2319, N299);
nand NAND2_2116 (N2347, N2319, N2112);
nand NAND2_2117 (N2348, N2330, N2300);
nand NAND2_2118 (N2349, N2331, N2301);
nand NAND2_2119 (N2350, N2332, N2302);
nand NAND2_2120 (N2351, N2333, N2303);
nand NAND2_2121 (N2352, N2335, N2304);
nand NAND2_2122 (N2353, N2337, N2305);
nand NAND2_2123 (N2354, N2339, N2306);
nand NAND2_2124 (N2355, N2341, N2307);
nand NAND2_2125 (N2356, N2343, N2308);
nand NAND2_2129 (N2371, N214,  N2360);
nand NAND2_2130 (N2372, N2360, N227);
nand NAND2_2131 (N2373, N2360, N240);
nand NAND2_2132 (N2374, N2360, N253);
nand NAND2_2133 (N2375, N2360, N266);
nand NAND2_2134 (N2376, N2360, N279);
nand NAND2_2135 (N2377, N2360, N292);
nand NAND2_2136 (N2378, N2360, N2105);
nand NAND2_2137 (N2379, N2360, N2115);
nand NAND3_2156 (N2428, N2399, N2393, N2419);
nand NAND4_2138 (N2380, N24,   N2242, N2334, N2371);
nand NAND4_2139 (N2381, N2246, N2336, N2372, N217);
nand NAND4_2140 (N2386, N2250, N2338, N2373, N230);
nand NAND4_2141 (N2393, N2254, N2340, N2374, N243);
nand NAND4_2142 (N2399, N2255, N2342, N2375, N256);
nand NAND4_2143 (N2404, N2256, N2344, N2376, N269);
nand NAND4_2144 (N2407, N2257, N2345, N2377, N282);
nand NAND4_2145 (N2411, N2258, N2346, N2378, N295);
nand NAND4_2146 (N2414, N2259, N2347, N2379, N2108);
nand NAND4_2155 (N2425, N2386, N2393, N2418, N2399);
nand NAND4_2157 (N2429, N2386, N2393, N2407, N2420);
nand NAND4_2158 (N2430, N2381, N2386, N2422, N2399);
nand NAND4_2159 (N2431, N2381, N2386, N2425, N2428);
nand NAND4_2160 (N2432, N2381, N2422, N2425, N2429);
and  AND8_2148  (N2416, N2381, N2386, N2393, N2399, N2404, N2407, N2411, N2414);
and  AND9_246   (N2199, N2154, N2159, N2162, N2165, N2168, N2171, N2174, N2177, N2180);
and  AND9_286   (N2296, N2260, N2264, N2267, N2270, N2273, N2276, N2279, N2282, N2285);
and  AND9_2126  (N2357, N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356);

endmodule
