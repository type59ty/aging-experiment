`timescale 1ns/10ps
//`include "c17.v"

`define cycle 10.0
`define terminate_cycle 400000//200000 // Modify your terminate ycle here

module c2670_testfixture;

`define in_file "c2670/rand_input_vector_c2670_0.out"
`define out_file "c2670/rand_output_vector_c2670_0.out"

parameter vec_width = 233;
parameter vec_length = 8;

reg clk = 0;


reg [vec_width-1:0] input_vec_mem [0:vec_length-1];
reg [vec_width-1:0] vec;


wire n398,n400,n401,n419,n420,n456,n457,n458,n487,n488,
     n489,n490,n491,n492,n493,n494,n792,n799,n805,n1026,
     n1028,n1029,n1269,n1277,n1448,n1726,n1816,n1817,n1818,n1819,
     n1820,n1821,n1969,n1970,n1971,n2010,n2012,n2014,n2016,n2018,
     n2020,n2022,n2387,n2388,n2389,n2390,n2496,n2643,n2644,n2891,
     n2925,n2970,n2971,n3038,n3079,n3546,n3671,n3803,n3804,n3809,
     n3851,n3875,n3881,n3882,n143_O,n144_O,n145_O,n146_O,n147_O,n148_O,
     n149_O,n150_O,n151_O,n152_O,n153_O,n154_O,n155_O,n156_O,n157_O,n158_O,
     n159_O,n160_O,n161_O,n162_O,n163_O,n164_O,n165_O,n166_O,n167_O,n168_O,
     n169_O,n170_O,n171_O,n172_O,n173_O,n174_O,n175_O,n176_O,n177_O,n178_O,
     n179_O,n180_O,n181_O,n182_O,n183_O,n184_O,n185_O,n186_O,n187_O,n188_O,
     n189_O,n190_O,n191_O,n192_O,n193_O,n194_O,n195_O,n196_O,n197_O,n198_O,
     n199_O,n200_O,n201_O,n202_O,n203_O,n204_O,n205_O,n206_O,n207_O,n208_O,
     n209_O,n210_O,n211_O,n212_O,n213_O,n214_O,n215_O,n216_O,n217_O,n218_O;

		 

initial begin
	//$timeformat(-9, 1, " ns", 9); //Display time in nanoseconds
	$readmemb(`in_file, input_vec_mem );
end

always #(`cycle/2) clk = ~clk;

c2670 c2670_1 (.N1(vec[232]),.N2(vec[231]),.N3(vec[230]),.N4(vec[229]),.N5(vec[228]),.N6(vec[227]),.N7(vec[226]),.N8(vec[225]),.N11(vec[224]),.N14(vec[223]),
              .N15(vec[222]),.N16(vec[221]),.N19(vec[220]),.N20(vec[219]),.N21(vec[218]),.N22(vec[217]),.N23(vec[216]),.N24(vec[215]),.N25(vec[214]),.N26(vec[213]),
              .N27(vec[212]),.N28(vec[211]),.N29(vec[210]),.N32(vec[209]),.N33(vec[208]),.N34(vec[207]),.N35(vec[206]),.N36(vec[205]),.N37(vec[204]),.N40(vec[203]),
              .N43(vec[202]),.N44(vec[201]),.N47(vec[200]),.N48(vec[199]),.N49(vec[198]),.N50(vec[197]),.N51(vec[196]),.N52(vec[195]),.N53(vec[194]),.N54(vec[193]),
              .N55(vec[192]),.N56(vec[191]),.N57(vec[190]),.N60(vec[189]),.N61(vec[188]),.N62(vec[187]),.N63(vec[186]),.N64(vec[185]),.N65(vec[184]),.N66(vec[183]),
              .N67(vec[182]),.N68(vec[181]),.N69(vec[180]),.N72(vec[179]),.N73(vec[178]),.N74(vec[177]),.N75(vec[176]),.N76(vec[175]),.N77(vec[174]),.N78(vec[173]),
              .N79(vec[172]),.N80(vec[171]),.N81(vec[170]),.N82(vec[169]),.N85(vec[168]),.N86(vec[167]),.N87(vec[166]),.N88(vec[165]),.N89(vec[164]),.N90(vec[163]),
              .N91(vec[162]),.N92(vec[161]),.N93(vec[160]),.N94(vec[159]),.N95(vec[158]),.N96(vec[157]),.N99(vec[156]),.N100(vec[155]),.N101(vec[154]),.N102(vec[153]),
              .N103(vec[152]),.N104(vec[151]),.N105(vec[150]),.N106(vec[149]),.N107(vec[148]),.N108(vec[147]),.N111(vec[146]),.N112(vec[145]),.N113(vec[144]),.N114(vec[143]),
              .N115(vec[142]),.N116(vec[141]),.N117(vec[140]),.N118(vec[139]),.N119(vec[138]),.N120(vec[137]),.N123(vec[136]),.N124(vec[135]),.N125(vec[134]),.N126(vec[133]),
              .N127(vec[132]),.N128(vec[131]),.N129(vec[130]),.N130(vec[129]),.N131(vec[128]),.N132(vec[127]),.N135(vec[126]),.N136(vec[125]),.N137(vec[124]),.N138(vec[123]),
              .N139(vec[122]),.N140(vec[121]),.N141(vec[120]),.N142(vec[119]),.N219(vec[118]),.N224(vec[117]),.N227(vec[116]),.N230(vec[115]),.N231(vec[114]),.N234(vec[113]),
              .N237(vec[112]),.N241(vec[111]),.N246(vec[110]),.N253(vec[109]),.N256(vec[108]),.N259(vec[107]),.N262(vec[106]),.N263(vec[105]),.N266(vec[104]),.N269(vec[103]),
              .N272(vec[102]),.N275(vec[101]),.N278(vec[100]),.N281(vec[99]),.N284(vec[98]),.N287(vec[97]),.N290(vec[96]),.N294(vec[95]),.N297(vec[94]),.N301(vec[93]),
              .N305(vec[92]),.N309(vec[91]),.N313(vec[90]),.N316(vec[89]),.N319(vec[88]),.N322(vec[87]),.N325(vec[86]),.N328(vec[85]),.N331(vec[84]),.N334(vec[83]),
              .N337(vec[82]),.N340(vec[81]),.N343(vec[80]),.N346(vec[79]),.N349(vec[78]),.N352(vec[77]),.N355(vec[76]),.N143_I(vec[75]),.N144_I(vec[74]),.N145_I(vec[73]),
              .N146_I(vec[72]),.N147_I(vec[71]),.N148_I(vec[70]),.N149_I(vec[69]),.N150_I(vec[68]),.N151_I(vec[67]),.N152_I(vec[66]),.N153_I(vec[65]),.N154_I(vec[64]),.N155_I(vec[63]),
              .N156_I(vec[62]),.N157_I(vec[61]),.N158_I(vec[60]),.N159_I(vec[59]),.N160_I(vec[58]),.N161_I(vec[57]),.N162_I(vec[56]),.N163_I(vec[55]),.N164_I(vec[54]),.N165_I(vec[53]),
              .N166_I(vec[52]),.N167_I(vec[51]),.N168_I(vec[50]),.N169_I(vec[49]),.N170_I(vec[48]),.N171_I(vec[47]),.N172_I(vec[46]),.N173_I(vec[45]),.N174_I(vec[44]),.N175_I(vec[43]),
              .N176_I(vec[42]),.N177_I(vec[41]),.N178_I(vec[40]),.N179_I(vec[39]),.N180_I(vec[38]),.N181_I(vec[37]),.N182_I(vec[36]),.N183_I(vec[35]),.N184_I(vec[34]),.N185_I(vec[33]),
              .N186_I(vec[32]),.N187_I(vec[31]),.N188_I(vec[30]),.N189_I(vec[29]),.N190_I(vec[28]),.N191_I(vec[27]),.N192_I(vec[26]),.N193_I(vec[25]),.N194_I(vec[24]),.N195_I(vec[23]),
              .N196_I(vec[22]),.N197_I(vec[21]),.N198_I(vec[20]),.N199_I(vec[19]),.N200_I(vec[18]),.N201_I(vec[17]),.N202_I(vec[16]),.N203_I(vec[15]),.N204_I(vec[14]),.N205_I(vec[13]),
              .N206_I(vec[12]),.N207_I(vec[11]),.N208_I(vec[10]),.N209_I(vec[9]),.N210_I(vec[8]),.N211_I(vec[7]),.N212_I(vec[6]),.N213_I(vec[5]),.N214_I(vec[4]),.N215_I(vec[3]),
              .N216_I(vec[2]),.N217_I(vec[1]),.N218_I(vec[0]),
							.N398(n398),.N400(n400),.N401(n401),.N419(n419),.N420(n420),.N456(n456),.N457(n457),
              .N458(n458),.N487(n487),.N488(n488),.N489(n489),.N490(n490),.N491(n491),.N492(n492),.N493(n493),.N494(n494),.N792(n792),
              .N799(n799),.N805(n805),.N1026(n1026),.N1028(n1028),.N1029(n1029),.N1269(n1269),.N1277(n1277),.N1448(n1448),.N1726(n1726),.N1816(n1816),
              .N1817(n1817),.N1818(n1818),.N1819(n1819),.N1820(n1820),.N1821(n1821),.N1969(n1969),.N1970(n1970),.N1971(n1971),.N2010(n2010),.N2012(n2012),
              .N2014(n2014),.N2016(n2016),.N2018(n2018),.N2020(n2020),.N2022(n2022),.N2387(n2387),.N2388(n2388),.N2389(n2389),.N2390(n2390),.N2496(n2496),
              .N2643(n2643),.N2644(n2644),.N2891(n2891),.N2925(n2925),.N2970(n2970),.N2971(n2971),.N3038(n3038),.N3079(n3079),.N3546(n3546),.N3671(n3671),
              .N3803(n3803),.N3804(n3804),.N3809(n3809),.N3851(n3851),.N3875(n3875),.N3881(n3881),.N3882(n3882),.N143_O(n143_O),.N144_O(n144_O),.N145_O(n145_O),
              .N146_O(n146_O),.N147_O(n147_O),.N148_O(n148_O),.N149_O(n149_O),.N150_O(n150_O),.N151_O(n151_O),.N152_O(n152_O),.N153_O(n153_O),.N154_O(n154_O),.N155_O(n155_O),
              .N156_O(n156_O),.N157_O(n157_O),.N158_O(n158_O),.N159_O(n159_O),.N160_O(n160_O),.N161_O(n161_O),.N162_O(n162_O),.N163_O(n163_O),.N164_O(n164_O),.N165_O(n165_O),
              .N166_O(n166_O),.N167_O(n167_O),.N168_O(n168_O),.N169_O(n169_O),.N170_O(n170_O),.N171_O(n171_O),.N172_O(n172_O),.N173_O(n173_O),.N174_O(n174_O),.N175_O(n175_O),
              .N176_O(n176_O),.N177_O(n177_O),.N178_O(n178_O),.N179_O(n179_O),.N180_O(n180_O),.N181_O(n181_O),.N182_O(n182_O),.N183_O(n183_O),.N184_O(n184_O),.N185_O(n185_O),
              .N186_O(n186_O),.N187_O(n187_O),.N188_O(n188_O),.N189_O(n189_O),.N190_O(n190_O),.N191_O(n191_O),.N192_O(n192_O),.N193_O(n193_O),.N194_O(n194_O),.N195_O(n195_O),
              .N196_O(n196_O),.N197_O(n197_O),.N198_O(n198_O),.N199_O(n199_O),.N200_O(n200_O),.N201_O(n201_O),.N202_O(n202_O),.N203_O(n203_O),.N204_O(n204_O),.N205_O(n205_O),
              .N206_O(n206_O),.N207_O(n207_O),.N208_O(n208_O),.N209_O(n209_O),.N210_O(n210_O),.N211_O(n211_O),.N212_O(n212_O),.N213_O(n213_O),.N214_O(n214_O),.N215_O(n215_O),
              .N216_O(n216_O),.N217_O(n217_O),.N218_O(n218_O) );							

integer i=0;
always @ (posedge clk) begin
	vec = input_vec_mem[i];
	$monitor(vec);
	i = i + 1;

end

always @ (negedge clk)begin
	$fdisplay ( fh_w, n398,n400,n401,n419,n420,n456,n457,n458,n487,n488,
	                  n489,n490,n491,n492,n493,n494,n792,n799,n805,n1026,
                    n1028,n1029,n1269,n1277,n1448,n1726,n1816,n1817,n1818,n1819,
                    n1820,n1821,n1969,n1970,n1971,n2010,n2012,n2014,n2016,n2018,
                    n2020,n2022,n2387,n2388,n2389,n2390,n2496,n2643,n2644,n2891,
                    n2925,n2970,n2971,n3038,n3079,n3546,n3671,n3803,n3804,n3809,
                    n3851,n3875,n3881,n3882,n143_O,n144_O,n145_O,n146_O,n147_O,n148_O,
                    n149_O,n150_O,n151_O,n152_O,n153_O,n154_O,n155_O,n156_O,n157_O,n158_O,
                    n159_O,n160_O,n161_O,n162_O,n163_O,n164_O,n165_O,n166_O,n167_O,n168_O,
                    n169_O,n170_O,n171_O,n172_O,n173_O,n174_O,n175_O,n176_O,n177_O,n178_O,
                    n179_O,n180_O,n181_O,n182_O,n183_O,n184_O,n185_O,n186_O,n187_O,n188_O,
                    n189_O,n190_O,n191_O,n192_O,n193_O,n194_O,n195_O,n196_O,n197_O,n198_O,
                    n199_O,n200_O,n201_O,n202_O,n203_O,n204_O,n205_O,n206_O,n207_O,n208_O,
                    n209_O,n210_O,n211_O,n212_O,n213_O,n214_O,n215_O,n216_O,n217_O,n218_O);	
	if(i == vec_length)begin
		$finish;
	end
end

integer fh_w;
initial begin
	fh_w = $fopen(`out_file, "w");
end
 
initial begin
	//$fsdbDumpfile("SET.fsdb");
	//$fsdbDumpvars;
	//$fsdbDumpMDA;
	$dumpfile("test_result.vcd");
    $dumpvars;

end
endmodule
